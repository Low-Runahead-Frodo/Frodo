module AddrLUT (
    input       [3:0]   index,
    output  reg [13:0]  addr
);
    always @(*) begin
        case (index)
            4'b0000: addr = 14'b00_0000_0000_0000;
            4'b0001: addr = 14'b00_0000_0000_0000;
            4'b0010: addr = 14'b01_0000_0100_0000;
            4'b0011: addr = 14'b11_0000_0000_0000;
            4'b0100: addr = 14'b00_0000_0000_0100;
            4'b0101: addr = 14'b00_0000_0000_0101;
            4'b0110: addr = 14'b00_0000_0000_0110;
            4'b0111: addr = 14'b00_0000_0000_0111;
            4'b1000: addr = 14'b00_0000_0000_1000;
            4'b1001: addr = 14'b00_0000_0000_1001;
            4'b1010: addr = 14'b00_0000_0000_1010;
            4'b1011: addr = 14'b00_0000_0000_1011;            
            4'b1100: addr = 14'b00_0000_0000_1100;            
            4'b1101: addr = 14'b00_0000_0000_1101;            
            4'b1110: addr = 14'b00_0000_0000_1110;              
            4'b1111: addr = 14'b11_0000_0110_0000;              
        endcase
    end
endmodule